library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity RCA_Input is

end RCA_Input;

architecture input of RCA_Input is

begin

end input;