library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity RCA_to_USB is

end RCA_to_USB;

architecture USB_convert of RCA_to_USB is

begin

end USB_convert;