library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity RCA_to_HDMI is

end RCA_to_HDMI;

architecture HDMI_convert of RCA_to_HDMI is

begin

end HDMI_convert;